`timescale 1ns / 1ps


module gp1(input wire a, b, output wire g, p);
    assign g = a & b; 
    assign p = a | b; 
endmodule

module gp4(input wire [3:0] gin, pin,
           input wire cin,
           output wire gout, pout,
           output wire [2:0] cout);

    wire [3:0] c_internal;
    assign c_internal[0] = cin;
    assign c_internal[1] = gin[0] | (pin[0] & c_internal[0]);
    assign c_internal[2] = gin[1] | (pin[1] & c_internal[1]);
    assign c_internal[3] = gin[2] | (pin[2] & c_internal[2]);

    assign cout[0] = c_internal[1];
    assign cout[1] = c_internal[2];
    assign cout[2] = c_internal[3];

    assign gout = gin[3] | (pin[3] & c_internal[3]);
    assign pout = pin[0] & pin[1] & pin[2] & pin[3];
endmodule

module gp8(input wire [7:0] gin, pin,
           input wire cin,
           output wire gout, pout,
           output wire [6:0] cout);

    wire [7:0] c_internal;
    assign c_internal[0] = cin;
    assign c_internal[1] = gin[0] | (pin[0] & c_internal[0]);
    // Corrected loop 
    genvar i;
    generate
        for (i = 1; i < 7; i = i + 1) begin : loop
            assign c_internal[i + 1] = gin[i] | (pin[i] & c_internal[i]);
        end
    endgenerate

    assign cout = c_internal[1:7]; // Correctly assign the internal carries to cout

    assign gout = gin[7] | (pin[7] & c_internal[7]);
    assign pout = &pin; // AND all propagate signals together
endmodule


module cla(input wire [31:0] a, b,
           input wire cin,
           output wire [31:0] sum);

    wire [31:0] g, p; // Generate and propagate for each bit
    wire [31:0] c; // Carry for each bit position, c[0] is cin
    wire [7:0] g8, p8; // Generate and propagate for 8-bit segments
    wire [3:0] cout8; // Carry out between 8-bit segments

    // Instantiate gp1 modules for each bit
    genvar i;
    generate
        for (i = 0; i < 32; i = i + 1) begin : gp1_gen
            gp1 gp1_inst(.a(a[i]), .b(b[i]), .g(g[i]), .p(p[i]));
        end
    endgenerate

    // Instantiate gp8 modules for each 8-bit segment
    gp8 gp8_inst0(.gin(g[7:0]), .pin(p[7:0]), .cin(cin), .gout(g8[0]), .pout(p8[0]), .cout(cout8[0]));
    gp8 gp8_inst1(.gin(g[15:8]), .pin(p[15:8]), .cin(cout8[0]), .gout(g8[1]), .pout(p8[1]), .cout(cout8[1]));
    gp8 gp8_inst2(.gin(g[23:16]), .pin(p[23:16]), .cin(cout8[1]), .gout(g8[2]), .pout(p8[2]), .cout(cout8[2]));
    gp8 gp8_inst3(.gin(g[31:24]), .pin(p[31:24]), .cin(cout8[2]), .gout(g8[3]), .pout(p8[3]), .cout(cout8[3]));

    // Calculate carry for the entire 32-bit operation, ensuring c[0] is cin
    assign c[0] = cin;
    
    // Intermediate carries within 8-bit segments should be properly calculated
    generate
        for (i = 1; i < 32; i = i + 1) begin : carry_gen
            if (i % 8 == 0) begin
                assign c[i] = cout8[i/8-1]; // Use cout8 from gp8 instances for carries at 8, 16, 24
            end else begin
                assign c[i] = g[i-1] | (p[i-1] & c[i-1]); // Calculate intermediate carries based on generate and propagate
            end
        end
    endgenerate

    // Calculate sum
    generate
        for (i = 0; i < 32; i = i + 1) begin : sum_gen
            assign sum[i] = a[i] ^ b[i] ^ c[i];
        end
    endgenerate

endmodule
